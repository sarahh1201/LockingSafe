library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity top is 
end top; 

architecture arch of top is 
end arch;